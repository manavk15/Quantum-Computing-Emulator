
                                               
`define Q_STATE_OUTPUT_SRAM_ADDRESS_UPPER_BOUND 32
`define Q_STATE_OUTPUT_SRAM_DATA_UPPER_BOUND  128
                                             
`define Q_STATE_INPUT_SRAM_ADDRESS_UPPER_BOUND 32
`define Q_STATE_INPUT_SRAM_DATA_UPPER_BOUND    128
                                             
`define SCRATCHPAD_SRAM_ADDRESS_UPPER_BOUND    32
`define SCRATCHPAD_SRAM_DATA_UPPER_BOUND       128
                                             
`define Q_GATES_SRAM_ADDRESS_UPPER_BOUND       32
`define Q_GATES_SRAM_DATA_UPPER_BOUND          128
